64x64y
9x37y
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111101111111111111111111111111111111
1111111111110001111111111000000000000110011111111111111111111111
1111111111000000000000000000000000000000000000011111111222001111
1111111100000000000000000000000000000000000000000111111200001111
1111111100000000000000000000000000000000000000000000111200001111
1111111000000000000000000000000000000000000000000000111200001111
1111110000000000000000000000000000000000000000000000111100001111
1111100000000000000000000000000000000000000000000000001110000111
1111100000000000011111111111111111111111111111000000000110000011
1111100000000000011111111111111111111111111111100000000000000011
1111100000000000011111111111111111111111111111000000000000000111
1111100000000000011111111111111111111111111000000000000000001111
1111000000000000011110011111111111111111111000000000000000001111
1111100000000000111110111111111111111111110000001000000000011111
1111000000000000111100000111111111111110000000001000000000011111
1111100000000000111100000111111111111000000000001100000000001111
1111000000000001111100000011111111110000000000001100000000000111
1111000000000001112200000011111111100000000000001110000000000111
1111000000000001112200000001111111000000000000000110000000001111
1110000000000001110000000001111100000000000000000100000000001111
1110000000000011110000000001111000000000000000000110000000001111
1111000000000011110000000001110000000000000000000110000000000111
1111000000000011100000000001110000000000000000000110000000000111
1111100000000111000000000001110000000000000000000110000000000111
1111000040000111000000000001100000000001000000000110000000000111
1111100000000111000000000001000000000011000000000110000000000111
1111110000001110000000000000000000000111000000000111000000000111
1111111111111110000000000000000000001111000000000111000000400111
1111111111101000000000000000000000001111000000000111000000000111
1111011000000000000000000000000000001111000000000110000000000111
1110000000000000000000000000000000001110000000000110000000000111
1111000000000000000100001000000000001110000000000111000000000111
1110000000000000000100101000000000001110000000000111000000000111
1110000000000000000101001100000000001110000000000111000000000111
1110000000000000000100101010000000011110000000000111000000000011
1110000000000000000000000000000000011110000000000111000000000011
1110000003000000000000000000000000011100000000000111000000000011
1111100000000000010000000000000000011110000000000111000000000111
1111100000000000111000000000000000011110000000000111000000000011
1111100000000011110000000000000000011110000000000111000000000011
1111000000000011110000000000000000111110000000000111000000000111
1111100000000111110000000000000000111110000000000111000000000111
1111110000111111111100000000000000111110000000000111000000000111
1111111000111111110000000000000000111111000000000111000000000111
1111111100011111111111111111000000111111000000000111000000000001
1111111111111111111111111111111100011111000000000111000000000011
1111111111111111111111111111111110111110000000000111000000000011
1111100000000000000000000001111111111110000000000111000000000011
1111100000000000000000000000111111111110000000000111000000000011
1111100000000000000000000000001111111100000000000011000000000011
1111000000000000000000000000000111111000000000000011000000000011
1111000000400000000000000000000000000000000000000010000000000011
1111110000000000000000000000000000000000000000000000000000000011
1111101000000000000000001000000000000000000000000000000000000011
1111100000000000111100000000000000000000000000000000000000000011
1111111000000001111110000000000000000000000000000000000000000011
1111110000000011111111000000000000000000000000011000000000000111
1111110000001111111111101000000000000000000001101111100000000111
1111111111111111111111111110000000000000000011111111111111111111
1111111111111111111111111220000110000000000111111111111111111111
1111111111111111111111111222001111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
