16x16y
2222222222222222
2111111211111112
2111111211111112
2111111211111112
2111111211111112
2112111211111112
2112111211111112
2112111211111112
2112111211111112
2112111211111112
2112111111111112
2112111111111112
2112111111111112
2112111111111112
2112111111111111
2222222222222222
