64x32y
2222222222222222222222222222222222222222222222222222222222222222
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111111211211111111111121121111111111112112111111111111
2222222222222222222222222222222222222222222222222222222222222222
2222222222222222222222222222222222222222222222222222222222222222
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111111211211111111111121121111111111112112111111111111
2222222222222222222222222222222222222222222222222222222222222222
