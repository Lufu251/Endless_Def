64x64y
2222211111111111111111111111111111111111111111111111111111111111
2111111111111111111111111111111111111111111111111111111111111111
2111121111111111111111111111111111111111111111111111111111111111
2111121111111111111111111111111111111111111111111111111111111111
2111121111111111111111111111111111111111111111111111111111111111
2111111111111111111111111111111111111111111111111111111111111111
2111121111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111
1111111111111111111111111111111111111111111111111111111111111111


32x32y
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111
11111111111111111111111111111111


128x64y
22222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111111111111211111112211111121111111111111112111111111111111211111111111111121111111221111112111111111111111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111112112111111111111111211111111111121121111111111112112111111111111211211111111111111121111111111112112111111111111
22222222222122222222222222122222222222222212222222222222122222222222222222212222222222222212222222222222221222222222222212222222
22222222222122222222222222122222222222222212222222222222122222222222222222212222222222222212222222222222221222222222222212222222
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111112112111111111111211211111111111121121111111111112112111111111111211211111111111121121111111111112112111111111111
22222222222122222222222222222222222222222212222222222222222222222222222222212222222222222222222222222222222122222222222222222222
22222222222222222222222222222222222222222212222222222222222222222222222222222222222222222222222222222222222122222222222222222222
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111111111111211111112211111121111111111111112111111111111111211111111111111121111111221111112111111111111111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111112112111111111111111211111111111121121111111111112112111111111111211211111111111111121111111111112112111111111111
22222222222122222222222222122222222222222212222222222222122222222222222222212222222222222212222222222222221222222222222212222222
22222222222122222222222222122222222222222212222222222222122222222222222222212222222222222212222222222222221222222222222212222222
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21111112111111122111111211111112211111121111111221111112111111122111111211111112211111121111111221111112111111122111111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121112111111122112111211111112211211121111111221121112111111122112111211111112211211121111111221121112111111122112111211111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111122112111111111112211211111111111221121111111111122112111111111112211211111111111221121111111111122112111111111112
21121111111111112112111111111111211211111111111121121111111111112112111111111111211211111111111121121111111111112112111111111111
22222222222122222222222222222222222222222222222222222222222222222222222222212222222222222222222222222222222222222222222222222222






64x32y
2222222222222222222222222222222222222222222222222222222222222222
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111111211211111111111121121111111111112112111111111111
2222222222222222222222222222222222222222222222222222222222222222
2222222222222222222222222222222222222222222222222222222222222222
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2111111211111112211111121111111221111112111111122111111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111211111112211211121111111221121112111111122112111211111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111112211211111111111221121111111111122112111111111112
2112111111111111211211111111111121121111111111112112111111111111
2222222222222222222222222222222222222222222222222222222222222222
